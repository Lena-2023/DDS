module note2dds_1st_gen(CLK, NOTE, ADDER);

input wire CLK;
input wire [7:0] NOTE;
output reg [31:0] ADDER;

initial begin
           ADDER <= 32'd0;
end

always @ (posedge CLK) begin
           case(NOTE)
8'd00: ADDER <= 32'd02;
8'd01: ADDER <= 32'd02;
8'd02: ADDER <= 32'd03;
8'd03: ADDER <= 32'd03;
8'd04: ADDER <= 32'd03;
8'd05: ADDER <= 32'd03;
8'd06: ADDER <= 32'd03;
8'd07: ADDER <= 32'd04;
8'd08: ADDER <= 32'd04;
8'd09: ADDER <= 32'd04;
8'd010: ADDER <= 32'd04;
8'd011: ADDER <= 32'd05;
8'd012: ADDER <= 32'd05;
8'd013: ADDER <= 32'd05;
8'd014: ADDER <= 32'd06;
8'd015: ADDER <= 32'd06;
8'd016: ADDER <= 32'd06;
8'd017: ADDER <= 32'd07;
8'd018: ADDER <= 32'd07;
8'd019: ADDER <= 32'd08;
8'd020: ADDER <= 32'd08;
8'd021: ADDER <= 32'd09;
8'd022: ADDER <= 32'd09;
8'd023: ADDER <= 32'd010;
8'd024: ADDER <= 32'd010;
8'd025: ADDER <= 32'd011;
8'd026: ADDER <= 32'd012;
8'd027: ADDER <= 32'd013;
8'd028: ADDER <= 32'd013;
8'd029: ADDER <= 32'd014;
8'd030: ADDER <= 32'd015;
8'd031: ADDER <= 32'd016;
8'd032: ADDER <= 32'd017;
8'd033: ADDER <= 32'd018;
8'd034: ADDER <= 32'd019;
8'd035: ADDER <= 32'd020;
8'd036: ADDER <= 32'd021;
8'd037: ADDER <= 32'd023;
8'd038: ADDER <= 32'd024;
8'd039: ADDER <= 32'd026;
8'd040: ADDER <= 32'd027;
8'd041: ADDER <= 32'd029;
8'd042: ADDER <= 32'd031;
8'd043: ADDER <= 32'd032;
8'd044: ADDER <= 32'd034;
8'd045: ADDER <= 32'd036;
8'd046: ADDER <= 32'd039;
8'd047: ADDER <= 32'd041;
8'd048: ADDER <= 32'd043;
8'd049: ADDER <= 32'd046;
8'd050: ADDER <= 32'd049;
8'd051: ADDER <= 32'd052;
8'd052: ADDER <= 32'd055;
8'd053: ADDER <= 32'd058;
8'd054: ADDER <= 32'd062;
8'd055: ADDER <= 32'd065;
8'd056: ADDER <= 32'd069;
8'd057: ADDER <= 32'd073;
8'd058: ADDER <= 32'd078;
8'd059: ADDER <= 32'd082;
8'd060: ADDER <= 32'd087;
8'd061: ADDER <= 32'd093;
8'd062: ADDER <= 32'd098;
8'd063: ADDER <= 32'd0104;
8'd064: ADDER <= 32'd0110;
8'd065: ADDER <= 32'd0117;
8'd066: ADDER <= 32'd0124;
8'd067: ADDER <= 32'd0131;
8'd068: ADDER <= 32'd0139;
8'd069: ADDER <= 32'd0147;
8'd070: ADDER <= 32'd0156;
8'd071: ADDER <= 32'd0165;
8'd072: ADDER <= 32'd0175;
8'd073: ADDER <= 32'd0186;
8'd074: ADDER <= 32'd0197;
8'd075: ADDER <= 32'd0208;
8'd076: ADDER <= 32'd0221;
8'd077: ADDER <= 32'd0234;
8'd078: ADDER <= 32'd0248;
8'd079: ADDER <= 32'd0263;
8'd080: ADDER <= 32'd0278;
8'd081: ADDER <= 32'd0295;
8'd082: ADDER <= 32'd0312;
8'd083: ADDER <= 32'd0331;
8'd084: ADDER <= 32'd0351;
8'd085: ADDER <= 32'd0372;
8'd086: ADDER <= 32'd0394;
8'd087: ADDER <= 32'd0417;
8'd088: ADDER <= 32'd0442;
8'd089: ADDER <= 32'd0468;
8'd090: ADDER <= 32'd0496;
8'd091: ADDER <= 32'd0526;
8'd092: ADDER <= 32'd0557;
8'd093: ADDER <= 32'd0590;
8'd094: ADDER <= 32'd0625;
8'd095: ADDER <= 32'd0662;
8'd096: ADDER <= 32'd0702;
8'd097: ADDER <= 32'd0744;
8'd098: ADDER <= 32'd0788;
8'd099: ADDER <= 32'd0835;
8'd0100: ADDER <= 32'd0884;
8'd0101: ADDER <= 32'd0937;
8'd0102: ADDER <= 32'd0993;
8'd0103: ADDER <= 32'd01052;
8'd0104: ADDER <= 32'd01114;
8'd0105: ADDER <= 32'd01181;
8'd0106: ADDER <= 32'd01251;
8'd0107: ADDER <= 32'd01325;
8'd0108: ADDER <= 32'd01404;
8'd0109: ADDER <= 32'd01488;
8'd0110: ADDER <= 32'd01576;
8'd0111: ADDER <= 32'd01670;
8'd0112: ADDER <= 32'd01769;
8'd0113: ADDER <= 32'd01874;
8'd0114: ADDER <= 32'd01986;
8'd0115: ADDER <= 32'd02104;
8'd0116: ADDER <= 32'd02229;
8'd0117: ADDER <= 32'd02362;
8'd0118: ADDER <= 32'd02502;
8'd0119: ADDER <= 32'd02651;
8'd0120: ADDER <= 32'd02809;
8'd0121: ADDER <= 32'd02976;
8'd0122: ADDER <= 32'd03153;
8'd0123: ADDER <= 32'd03340;
8'd0124: ADDER <= 32'd03539;
8'd0125: ADDER <= 32'd03749;
8'd0126: ADDER <= 32'd03972;
8'd0127: ADDER <= 32'd04209;
8'd0128: ADDER <= 32'd04459;
8'd0129: ADDER <= 32'd04724;
8'd0130: ADDER <= 32'd05005;
8'd0131: ADDER <= 32'd05303;
8'd0132: ADDER <= 32'd05618;
8'd0133: ADDER <= 32'd05952;
8'd0134: ADDER <= 32'd06306;
8'd0135: ADDER <= 32'd06681;
8'd0136: ADDER <= 32'd07078;
8'd0137: ADDER <= 32'd07499;
8'd0138: ADDER <= 32'd07945;
8'd0139: ADDER <= 32'd08418;
8'd0140: ADDER <= 32'd08918;
8'd0141: ADDER <= 32'd09448;
8'd0142: ADDER <= 32'd010010;
8'd0143: ADDER <= 32'd010606;
8'd0144: ADDER <= 32'd011236;
8'd0145: ADDER <= 32'd011904;
8'd0146: ADDER <= 32'd012612;
8'd0147: ADDER <= 32'd013362;
8'd0148: ADDER <= 32'd014157;
8'd0149: ADDER <= 32'd014999;
8'd0150: ADDER <= 32'd015891;
8'd0151: ADDER <= 32'd016836;
8'd0152: ADDER <= 32'd017837;
8'd0153: ADDER <= 32'd018897;
8'd0154: ADDER <= 32'd020021;
8'd0155: ADDER <= 32'd021212;
8'd0156: ADDER <= 32'd022473;
8'd0157: ADDER <= 32'd023809;
8'd0158: ADDER <= 32'd025225;
8'd0159: ADDER <= 32'd026725;
8'd0160: ADDER <= 32'd028314;
8'd0161: ADDER <= 32'd029998;
8'd0162: ADDER <= 32'd031782;
8'd0163: ADDER <= 32'd033672;
8'd0164: ADDER <= 32'd035674;
8'd0165: ADDER <= 32'd037795;
8'd0166: ADDER <= 32'd040043;
8'd0167: ADDER <= 32'd042424;
           endcase
end

endmodule


module DDS( 
input wire CLK,
input wire RESET,
input wire [31:0] ADDER, 
output reg [31:0]  DDS 
);

always @ (posedge CLK or posedge RESET) begin
  if(RESET)
   DDS <= 0;
  else
   DDS <= DDS + ADDER;
end

endmodule


module TOP (
input wire CLK,
input wire RESET,

input wire [7:0] NOTE,
output wire [31:0] DDS 
);


    note2dds_1st_gen N2D (.CLK(CLK), .NOTE(NOTE), .ADDER(ADDER));
    DDS DDS1 (.CLK(CLK), .RESET(RESET), .ADDER(ADDER), .DDS(DDS));

endmodule
